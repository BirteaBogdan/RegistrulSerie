library verilog;
use verilog.vl_types.all;
entity test_sreg is
end test_sreg;
